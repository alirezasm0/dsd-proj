// Copyright (c) 2018  LulinChen, All Rights Reserved
// AUTHOR : 	LulinChen
// AUTHOR'S EMAIL : lulinchen@aliyun.com 
// Release history
// VERSION Date AUTHOR DESCRIPTION

`include "global.sv"

`define	MAX_PATH			256
module tb();

	parameter  FRAME_WIDTH = 112;
	parameter  FRAME_HEIGHT = 48;
	parameter  SIM_FRAMES = 2;
	reg						rstn;
	reg						clk;
	reg						ee_clk;
	
	wire		rstn_ee = rstn;
	initial begin
		rstn = `RESET_ACTIVE;
		#(`RESET_DELAY); 
		$display("T%d rstn done#############################", $time);
		rstn = `RESET_IDLE;
	end
	
	initial begin
		clk = 1;
		forever begin
			clk = ~clk;
			#(`CLK_PERIOD_DIV2);
		end
	end
	
	initial begin
		ee_clk = 1;
		forever begin
			ee_clk = ~ee_clk;
			#(`EE_CLOCK_PERIOD_DIV2);
		end
	end
	
	
	
	reg			[15:0]			frame_width_0;
	reg			[15:0]			frame_height_0;
	reg			[31:0]			pic_to_sim;
	reg		[`MAX_PATH*8-1:0]	sequence_name_0;

	
		
	itf_data_punch itf(clk);
	wire									go =  itf.go;
	wire									en =  itf.en;
	wire									first_data =  itf.first_data;
	wire									last_data =  itf.last_data;
	wire	[`WDP*`INPUT_NUM-1:0]			data_i =  itf.data_i;
	wire	[`WDP*`OUTPUT_NUM*`INPUT_NUM-1:0]			weight =  itf.weight;
	wire	[`WDP*`OUTPUT_NUM-1:0]							bias =  itf.bias;

	initial begin
		#(`RESET_DELAY)
		#(`RESET_DELAY)
		itf.drive_a_frame();
		#(`RESET_DELAY)
		itf.drive_a_frame();
		#(30000* `TIME_COEFF)
		$finish();
	end	
	

	conv #(
		.INPUT_NUM		(1),
		.OUTPUT_NUM		(`OUTPUT_NUM)
		)conv(
		.clk			(clk),
		.rstn			(rstn),
		.go				(go),
		.en				(en),
		.first_data		(first_data),
		.last_data		(last_data),
		.data_i			(data_i),
		.bias			(bias),
		.weight			(weight),
		.q              ()
		);
	
		
`ifdef DUMP_FSDB 
	initial begin
	$fsdbDumpfile("fsdb/xx.fsdb");
	$fsdbDumpvars();
	end
`endif
	
endmodule


interface itf_data_punch(input clk);
	logic									go;
	logic									en;
	logic									first_data;
	logic									last_data;
	logic	[0:`INPUT_NUM-1][`WD:0]			data_i;
	logic	[0:`OUTPUT_NUM-1][`WD:0]		weight;
	logic	[0:`OUTPUT_NUM-1][`WD:0]		bias;
	
	clocking cb@( `CLK_EDGE);
		output	go;
		output	en;
		output	first_data;
		output	last_data;
		output	data_i;
		output	weight;
		output	bias;
	endclocking	
	
	//task drive_a_frame(int INPUT_NUM, int OUTPUT_NUM);
	task drive_a_frame();
		
		logic [0:4][0:4][0:5][31:0] weight0 = {
   3,    49,    -2,    -2,    37,    42,  
 -28,   -19,   -36,    51,    20,     0,  
 -28,   -62,   -50,    -4,    70,    22,  
  20,   -36,    38,   -26,    68,   -43,  
 -13,    39,    18,   -47,    49,   -48,  

  19,    61,   -23,    17,   -45,    54,  
  37,   -45,   -29,    41,   -19,    29,  
   6,   -64,    13,   -24,   -58,   -20,  
   6,    -1,    -8,   -62,    34,   -38,  
  13,    61,    44,   -57,    28,   -56,  

  33,     3,    32,    -8,   -26,    50,  
  22,   -14,    -4,    -9,    -9,    62,  
  53,   -74,     7,    15,  -118,     6,  
  59,     8,    23,    -7,   -79,    45,  
  10,    25,    38,   -25,   -35,   -22,  

  40,     6,    46,   -16,    -6,    -6,  
  16,   -37,    53,    44,    14,     4,  
  75,   -32,    44,    63,   -36,     5,  
  29,    -4,    48,    43,   -14,   -20,  
   2,    21,    59,     0,   -40,    -1,  

  11,    -3,    22,    38,   -14,    43,  
  22,   -31,     0,    35,    15,     7,  
  34,   -44,     0,    39,    65,    63,  
  -1,    15,    26,    34,    -5,   -12,  
 -22,    19,    15,    19,     0,   -23  
		};
		
		logic [0:31][0:31][31:0] test	 = {
			   0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0, 
			   0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0, 
			   0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0, 
			   0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0, 
			   0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0, 
			   0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0, 
			   0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0, 
			   0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0, 
			   0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0, 
			   0,    0,    0,    0,    0,    0,    0,    0,   84,  185,  159,  151,   60,   36,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0, 
			   0,    0,    0,    0,    0,    0,    0,    0,  222,  254,  254,  254,  254,  241,  198,  198,  198,  198,  198,  198,  198,  198,  170,   52,    0,    0,    0,    0,    0,    0,    0,    0, 
			   0,    0,    0,    0,    0,    0,    0,    0,   67,  114,   72,  114,  163,  227,  254,  225,  254,  254,  254,  250,  229,  254,  254,  140,    0,    0,    0,    0,    0,    0,    0,    0, 
			   0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,   17,   66,   14,   67,   67,   67,   59,   21,  236,  254,  106,    0,    0,    0,    0,    0,    0,    0,    0, 
			   0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,   83,  253,  209,   18,    0,    0,    0,    0,    0,    0,    0,    0, 
			   0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,   22,  233,  256,   83,    0,    0,    0,    0,    0,    0,    0,    0,    0, 
			   0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,  129,  254,  238,   44,    0,    0,    0,    0,    0,    0,    0,    0,    0, 
			   0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,   59,  249,  254,   62,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0, 
			   0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,  133,  254,  187,    5,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0, 
			   0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    9,  205,  248,   58,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0, 
			   0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,  126,  254,  182,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0, 
			   0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,   75,  251,  240,   57,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0, 
			   0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,   19,  221,  254,  166,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0, 
			   0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    3,  203,  254,  219,   35,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0, 
			   0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,   38,  254,  254,   77,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0, 
			   0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,   31,  224,  254,  115,    1,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0, 
			   0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,  133,  254,  254,   52,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0, 
			   0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,   61,  242,  254,  254,   52,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0, 
			   0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,  121,  254,  254,  219,   40,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0, 
			   0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,  121,  254,  207,   18,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0, 
			   0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0, 
			   0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0, 
			   0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0,    0
		};
		
			//    kernel_w  kernel_h output_num  input_num
			logic [0:4][0:4][0:15][0:5][31:0] weight1 = {
				  29,    29,    39,     6,   -15,     0,  
				   8,     4,    -9,   -14,   -24,     4,  
				  27,   -22,   -35,    26,    -9,    23,  
				  28,   -26,    35,   -26,   -70,   -10,  
				 -31,    41,   -12,   -31,   -23,   -27,  
				  13,    34,    -7,    -8,   -12,   -26,  
				 -37,   -12,    22,     8,    40,   -12,  
				 -45,   -62,   -57,    18,    62,    14,  
				   0,     9,   -10,   -21,   -48,   -15,  
				  18,   -29,   -39,    15,    14,    12,  
				 -11,    -1,   -10,    20,    21,    24,  
				  -6,   -54,   -38,    22,    33,   -31,  
				  12,    21,   -14,   -20,     9,   -23,  
				  -1,    74,    13,     6,   -35,   -15,  
				   2,    58,   -29,   -58,    31,   -23,  
				  15,    26,    -6,     1,    -9,   -24,  

				 -24,    15,   -24,    47,   -11,    -3,  
				  18,    69,    -7,    -6,   -31,    -6,  
				 -66,     4,    27,    -7,   -22,    41,  
				  21,   -27,    53,     2,   -14,   -19,  
				  46,   -31,    22,    39,     7,     2,  
				 -36,    31,    -2,    11,    -7,   -40,  
				 -35,   -22,    29,     0,   -39,    35,  
				 -19,     0,   -25,    15,    63,   -19,  
				  23,   -24,   -10,     0,    36,    27,  
				 -38,   -48,    30,    -3,    26,    21,  
				 -26,    75,    -4,    -2,   -34,     8,  
				 -32,   -35,   -58,    13,   -16,   -11,  
				 -11,     8,   -15,    34,   -13,    12,  
				 -13,     9,   -41,   -35,    15,    23,  
				  27,    13,    18,    21,     4,   -12,  
				  27,    38,   -15,     0,     2,    -5,  

				 -28,     7,   -14,   -29,    -4,    -3,  
				 -27,    50,   -34,   -32,   -78,   -26,  
				  -2,    58,    26,   -11,   -36,   -21,  
				   0,   -13,     3,    41,   -14,    39,  
				   3,    -6,    19,    32,   -11,    50,  
				   0,    76,     0,    18,   -30,     2,  
				 -18,    10,   -11,     7,   -54,    -3,  
				 -14,    -6,   -49,   -44,    62,   -26,  
				   7,   -24,   -35,    41,    36,   -10,  
				  50,   -24,    23,    19,   -40,   -27,  
				  21,    38,    46,    22,   -34,   -11,  
				  -1,    -7,    -6,    13,    -8,   -38,  
				  18,   -66,     0,     5,    28,    38,  
				   8,    49,    28,   -23,    -8,   -39,  
				  20,   -13,   -30,   -27,    28,    35,  
				  28,   -55,    16,    47,   -13,    27,  

				 -32,     3,    -1,   -50,   -15,     0,  
				 -20,    -1,    33,   -14,  -109,   -37,  
				  16,    -1,   -22,    33,   -38,    48,  
				  24,    17,    32,    -6,   -39,   -23,  
				  17,   -10,    46,    -6,     8,    28,  
				  11,    52,   -28,   -25,    13,    45,  
				 -29,   -20,    -2,    23,   -45,     3,  
				 -34,     4,   -29,    -8,    48,   -22,  
				  11,    26,    24,     4,    66,   -27,  
				   8,   -22,    21,    10,   -15,     0,  
				 -19,    19,    -4,    12,   -63,   -11,  
				  21,    33,   -37,    27,    -5,    13,  
				  10,    -2,    10,    -7,   -31,    17,  
				  -6,    12,    33,    26,   -13,    -2,  
				  43,    -1,    30,    -1,    48,    12,  
				  -3,   -33,    42,    35,     0,    39,  

				  34,   -27,    -3,    10,   -27,    11,  
				  18,    11,    30,   -53,   -63,   -26,  
				   7,    55,    43,   -11,   -34,    24,  
				 -30,   -28,    33,    27,   -28,    -5,  
				  15,    -4,    28,     6,    26,    28,  
				   6,    63,   -48,    17,    54,   -39,  
				   4,     1,    -9,   -19,   -41,    -5,  
				 -50,   -31,     8,    -6,    15,   -34,  
				 -49,   -17,   -17,   -39,    34,   -28,  
				  20,   -31,     7,    15,   -49,    25,  
				  21,    18,    -6,    43,    21,   -27,  
				  18,    -2,     1,   -40,    12,     7,  
				 -45,   -10,   -58,     9,    -2,     7,  
				   7,    -4,    17,    10,    -8,    31,  
				  44,   -25,    38,    22,    15,     4,  
				  18,   -57,   -17,    35,   -23,    23,  


				  24,    33,    44,   -12,   -39,    -5,  
				  14,    19,   -20,   -44,   -41,   -16,  
				  -9,     8,   -46,   -25,   -37,    21,  
				  51,     0,   -15,    -4,     5,    14,  
				 -10,    -5,   -32,    38,     1,    31,  
				  15,   -29,   -19,   -13,    -5,   -34,  
				  28,   -23,    30,     5,   -10,    11,  
				  32,   -83,    47,    37,    60,    20,  
				   5,   -61,   -39,    50,   -14,    10,  
				 -22,    13,    44,    37,   -28,    -4,  
				   6,    -5,   -26,    41,    21,    19,  
				  25,   -57,    48,    -5,    13,   -26,  
				  -9,     0,   -24,    -4,    22,   -36,  
				  17,    10,    12,    60,    -8,    24,  
				   0,    12,    18,   -19,     2,   -30,  
				 -14,   -23,    17,    12,     2,    51,  

				   5,    46,    -8,    25,    11,     0,  
				  13,    74,   -16,   -25,  -114,   -41,  
				 -61,     5,    -5,    -3,   -31,    27,  
				  63,     2,     2,     1,    -6,    10,  
				  56,   -23,   -10,    25,   -49,    10,  
				 -35,    11,    -4,   -39,   -24,    18,  
				  48,     0,     0,   -50,     0,   -50,  
				 -28,   -67,    25,    -1,    37,     9,  
				 -45,   -71,   -40,     4,    65,   -26,  
				  18,   -17,     2,    11,     9,   -28,  
				 -14,   -36,    20,     6,    19,    -6,  
				   5,   -13,    34,    15,    13,   -11,  
				  10,    -1,     5,     4,    12,    -4,  
				  36,    -6,    39,    33,    13,     3,  
				 -24,    59,   -11,   -44,    56,   -32,  
				 -11,    26,    -6,   -29,     7,   -22,  

				 -22,     2,    36,   -14,    12,   -25,  
				 -18,    51,     0,   -25,  -114,    -2,  
				  37,     7,     0,   -24,    -1,   -26,  
				   5,   -26,     9,   -23,    15,    33,  
				  -1,   -14,    17,   -12,   -49,    25,  
				 -27,    37,    14,   -19,    14,     4,  
				  -6,   -28,    16,   -35,   -22,     2,  
				  13,   -41,    16,    18,     1,   -31,  
				 -12,   -37,   -11,    30,    47,    27,  
				   9,     3,    10,    11,     2,    30,  
				 -53,    30,    20,   -56,   -29,     3,  
				  -3,   -28,    32,    34,   -15,    16,  
				   2,   -10,    31,    22,   -52,   -22,  
				  -2,   -39,   -16,    28,   -17,    19,  
				 -15,   -17,   -13,   -34,    48,   -39,  
				  15,    15,    10,     7,   -38,     3,  

				  11,    49,    33,   -67,   -42,   -61,  
				 -13,    77,   -14,   -33,   -44,    12,  
				  17,    -8,   -11,    21,    -4,     6,  
				   5,   -29,    35,    31,    38,    30,  
				  19,     0,   -14,    -8,     6,    27,  
				  16,    59,   -25,     9,   -29,    -2,  
				  45,   -34,    17,     6,    -5,     0,  
				  14,    -7,    14,    55,   -33,   -51,  
				 -13,   -67,   -17,     6,    95,    26,  
				 -21,   -26,    -5,    61,   -34,   -42,  
				   9,    12,     7,     5,   -37,    16,  
				  24,    -9,    -5,   -43,   -26,   -12,  
				  18,   -11,    10,    19,    16,    59,  
				  19,   -13,    -2,    16,   -21,   -18,  
				 -39,   -22,   -21,   -23,    40,   -11,  
				   3,     8,   -16,    55,   -14,     7,  

				  15,    -6,    26,   -14,   -64,    -9,  
				 -29,    68,   -26,     9,   -57,    48,  
				  28,    32,   -23,    48,   -19,    40,  
				  51,   -12,   -24,   -10,    30,    21,  
				  26,    -7,    -9,    29,     2,    22,  
				 -42,    59,   -43,   -29,    -9,    -8,  
				 -22,   -26,    32,    -4,    35,    20,  
				 -20,   -20,    -4,     1,    -6,    19,  
				 -36,   -45,   -56,   -47,    48,    -4,  
				  -9,    34,    21,    44,   -17,    16,  
				   2,     0,    -9,    67,   -10,    56,  
				  13,     5,   -15,   -42,    29,    -2,  
				 -22,    -8,   -39,    38,    50,    18,  
				  57,   -12,     7,    37,    27,    13,  
				 -35,    49,    42,   -19,     3,   -29,  
				  43,     1,    29,    19,   -52,    -5,  


				  -5,    31,   -14,    -8,    -5,    34,  
				 -19,    13,    -9,    13,   -75,    21,  
				 -35,    31,    12,   -45,    -6,     9,  
				  13,   -11,   -21,   -25,    88,   -10,  
				 -14,    -8,   -21,   -11,    36,   -40,  
				  16,    -7,     9,     0,    -3,    16,  
				  46,    21,    43,    -1,    -3,   -52,  
				  47,   -37,    21,    18,    13,   -27,  
				  -5,    -7,   -18,    26,    19,    19,  
				  36,   -18,   -20,     0,     4,    -1,  
				 -13,    18,   -15,   -17,    24,     3,  
				  18,   -13,     1,   -11,     0,   -28,  
				 -10,    -9,    24,    18,    23,   -43,  
				  15,   -12,    47,   -28,     7,   -10,  
				 -24,    10,   -10,   -19,   -14,    -3,  
				 -16,     4,   -24,     3,    22,    39,  

				 -12,   -22,   -14,   -23,   -23,    34,  
				 -13,    29,    20,    57,   -61,   -18,  
				  -6,    -8,    66,   -37,   -55,   -22,  
				   2,   -14,   -45,   -20,    47,   -22,  
				   2,    -2,   -37,   -69,    30,   -46,  
				 -15,   -39,   -27,   -14,     1,    -5,  
				  -4,     0,   -21,   -38,   -50,   -24,  
				  46,   -32,     8,   -15,    39,    41,  
				 -50,   -58,     8,    11,    42,   -37,  
				   9,   -41,    22,   -35,     7,    -4,  
				  14,    14,    12,    11,     2,   -54,  
				 -22,    -9,     4,   -34,    18,   -29,  
				  13,   -16,    18,   -11,    -1,   -24,  
				  15,    33,    31,    14,     3,     9,  
				   9,   -56,   -25,    31,     3,   -36,  
				  -2,     9,    -6,    -4,   -17,   -45,  

				  21,    28,    10,     2,   -25,   -48,  
				 -11,    23,    15,    59,   -18,   -10,  
				  18,     6,    31,     3,   -37,    31,  
				   3,   -19,   -33,    -9,    95,   -40,  
				 -46,     5,     3,   -13,     0,   -46,  
				 -15,    43,    -4,     0,    50,     8,  
				  -1,    -3,    15,    19,   -27,    33,  
				  11,   -30,     0,     6,    11,     0,  
				  -1,   -54,    -5,   -26,    53,    -4,  
				  16,   -38,    10,    43,    14,    27,  
				 -16,    33,    35,   -46,   -25,     8,  
				  -3,   -18,    38,     0,     0,    18,  
				  -8,    -5,    24,     0,    -1,   -21,  
				  21,    23,    27,   -16,     3,   -38,  
				   8,     9,   -40,   -13,    10,   -10,  
				  36,    -2,   -20,   -44,    12,    11,  

				  -8,    55,    10,   -14,   -45,     1,  
				  10,   -22,    10,    47,   -16,    42,  
				  23,    15,    32,    28,   -15,    17,  
				 -45,    -7,   -29,   -30,    29,    -9,  
				   5,    14,    30,     7,   -62,    26,  
				 -39,    22,   -18,   -47,     2,    -1,  
				  38,    55,     3,    -3,   -38,    12,  
				  44,   -21,     3,   -10,    -4,    -2,  
				  -7,   -17,    -2,    20,    53,     4,  
				   0,   -73,    21,    35,    17,   -11,  
				 -22,    35,     8,    42,   -53,   -15,  
				 -12,   -22,    -2,    -1,    15,    -2,  
				  -5,   -12,    26,    33,   -27,    10,  
				  14,   -13,     0,   -47,    -7,   -34,  
				 -49,   -10,   -15,     4,    34,    -8,  
				   7,    23,   -15,     6,    33,    -6,  

				  50,    69,    28,    -4,   -55,    36,  
				 -12,   -27,    47,    35,    11,    41,  
				 -47,    48,   -17,   -16,     1,    13,  
				  -5,    43,   -23,    -5,    65,    31,  
				  39,   -20,   -25,   -16,    -5,     9,  
				 -36,    -3,     7,    12,   -16,   -20,  
				   0,     0,   -36,     2,    27,   -27,  
				  40,   -16,    22,   -30,    54,   -15,  
				  41,   -23,    40,    49,    12,    -7,  
				  10,   -49,    12,     2,    19,    49,  
				   7,   -41,    15,     7,    -6,    45,  
				 -40,    -3,    18,    -6,   -23,     0,  
				   9,   -34,     6,     6,    24,    55,  
				 -15,    19,   -26,    20,     5,    20,  
				  29,    37,    -1,   -11,     5,    13,  
				  17,    31,    12,     9,   -42,    45,  


				   0,    55,   -44,     3,   -31,    51,  
				  -7,   -58,    35,    20,    -1,    29,  
				 -34,    14,    14,    17,   -36,    -7,  
				 -35,     8,   -49,   -23,    20,    -1,  
				 -64,   -65,   -25,   -29,     4,   -50,  
				  34,    -9,    -8,    35,   -62,   -16,  
				  -8,   -10,    39,    -8,   -39,   -31,  
				 -32,    47,   -13,    11,    15,   -49,  
				   5,   -71,    -1,    42,    13,    19,  
				  31,    -5,   -10,   -21,    19,    -1,  
				 -25,    -5,    37,   -18,     9,   -30,  
				  -1,   -23,   -18,    13,    85,    17,  
				  42,   -54,   -10,    31,   -45,   -57,  
				 -48,    -2,     5,   -37,    67,   -15,  
				  44,    11,    38,   -11,    -5,    16,  
				  19,    10,   -15,   -17,    60,   -28,  

				 -35,   -34,   -12,    -6,    13,    17,  
				  18,   -46,    39,    48,    40,    26,  
				  28,   -36,    48,   -14,  -107,    -9,  
				 -12,     0,   -35,    -4,    51,   -42,  
				 -57,     5,   -30,   -20,   -56,   -17,  
				   6,   -26,    13,     6,    28,    44,  
				  14,    30,    48,   -22,   -20,    16,  
				  17,   -16,    -2,    15,    -1,    -5,  
				  33,   -13,    15,    47,   -29,    55,  
				   0,   -25,     4,    24,    92,   -25,  
				   5,   -17,   -49,   -39,   -32,   -13,  
				  21,   -19,   -47,    29,    10,    14,  
				  -2,     2,    18,    -3,   -16,    -8,  
				 -49,    25,     5,   -35,    71,    11,  
				  22,   -39,    20,   -23,    22,    -9,  
				  -7,    34,   -31,    -9,   -23,    -9,  

				   2,     0,    -2,    -1,   -41,   -35,  
				 -21,   -28,     2,    42,    40,   -17,  
				  -7,    13,    55,   -24,   -45,     5,  
				 -27,   -13,   -12,     9,    27,   -66,  
				  -7,    27,    22,   -11,   -22,   -40,  
				   1,   -29,    34,    56,   -34,    -8,  
				  12,    48,    26,    -8,   -12,    45,  
				  57,     6,     9,    50,    16,    33,  
				  -6,   -14,    -5,   -44,   -15,    11,  
				   5,   -16,   -42,   -65,    42,    12,  
				 -25,    32,    16,     6,     3,   -28,  
				 -33,     4,   -20,    11,    67,    23,  
				   4,    -6,   -24,    -6,     7,   -14,  
				 -12,    14,   -23,    13,   -25,   -20,  
				 -38,   -35,   -19,    18,    15,   -32,  
				  15,    35,    18,   -57,   -47,   -44,  

				  18,    71,   -10,   -12,   -78,   -38,  
				  26,    -2,   -15,    21,    21,    26,  
				  -4,    65,   -51,    22,    -9,    39,  
				 -22,    -1,   -17,   -46,    35,   -50,  
				  33,    18,     3,    24,   -36,    55,  
				  -2,    15,    -3,    26,    14,   -17,  
				  -5,    60,   -17,     0,   -18,    42,  
				 -11,   -20,     3,   -31,    63,    13,  
				   9,   -16,    -9,    36,    29,    20,  
				  -5,     8,    43,   -34,    43,   -23,  
				 -47,     0,    13,   -48,     1,    -2,  
				  35,   -32,    30,    13,    -5,    29,  
				 -38,   -18,     3,   -43,    70,    -3,  
				 -67,    48,   -13,    17,     7,     0,  
				  -6,    30,    49,    -7,   -66,   -65,  
				  28,    20,    52,   -16,   -45,   -29,  

				  -1,    55,     4,    58,   -37,    48,  
				  34,   -19,     9,    48,    26,    -6,  
				 -29,    41,   -67,   -13,     5,    19,  
				 -29,    -1,   -18,    -3,   -36,   -19,  
				  16,    17,     0,     6,     6,    18,  
				  16,   -19,    51,     6,     0,    23,  
				   3,    22,    -2,    21,     3,   -17,  
				 -33,   -65,    15,    -4,    -2,    11,  
				  32,   -14,   -10,    33,     1,     0,  
				  24,   -18,    27,    13,    63,    15,  
				 -15,   -56,     4,    -2,   -20,   -12,  
				  22,    -9,    57,    25,   -61,   -28,  
				   0,   -34,   -17,    48,    -8,     9,  
				   7,    28,   -20,    -6,   -38,     0,  
				   7,    53,    54,   -25,   -91,   -44,  
				 -20,    49,   -28,    -6,   -14,    27,  


				  -9,    -3,   -15,   -17,    34,    -6,  
				  43,     2,   -12,   -16,    52,   -47,  
				  63,    14,     6,   -23,   -14,   -34,  
				  11,     5,   -10,   -26,   -39,     8,  
				  -8,     2,   -45,    -2,   -48,   -17,  
				   9,   -43,    18,   -32,    -5,   -21,  
				  13,     0,    42,     7,   -46,   -53,  
				   0,     1,   -35,    27,     6,     2,  
				 -23,    16,    25,    59,    54,    27,  
				 -19,   -53,   -46,   -13,   -10,   -35,  
				  37,    -5,    11,     4,   -12,   -10,  
				 -50,   -41,    12,    25,    51,    21,  
				   5,   -45,   -19,   -34,    45,    33,  
				 -15,   -15,   -29,    -5,    -4,    17,  
				  30,     3,   -38,   -21,    37,   -28,  
				  24,   -54,   -22,    37,    24,   -13,  

				 -27,   -21,   -33,   -21,   -29,   -19,  
				 -45,   -28,   -20,   -42,    34,     9,  
				  43,    16,   -26,   -11,   -17,    -9,  
				  33,    -8,     3,     0,   -41,    26,  
				 -11,   -34,    16,   -22,    22,   -16,  
				  17,   -32,   -10,    12,   -13,    39,  
				 -11,    57,     8,    11,   -29,    45,  
				  -2,    22,   -24,     4,    28,   -61,  
				  30,    40,    21,    14,     4,    60,  
				 -22,   -33,   -31,    32,    32,    -9,  
				 -20,   -29,    11,    -3,     0,    -6,  
				  24,   -29,    15,    28,    -1,   -31,  
				 -31,   -25,     6,    50,    47,   -10,  
				   0,   -36,   -21,   -41,    45,   -18,  
				  21,    20,   -49,    26,   -11,    22,  
				 -12,    -8,     3,     0,    21,   -21,  

				 -43,     6,   -34,    -3,    -6,   -14,  
				 -12,   -65,   -24,   -48,    79,    17,  
				   1,    43,   -45,    22,   -23,    12,  
				  16,   -36,    43,   -36,   -44,   -20,  
				  34,    30,    33,   -28,   -14,    -3,  
				  44,   -63,    36,    -8,   -13,    -1,  
				 -22,    43,   -24,   -16,   -26,   -23,  
				 -10,   -29,    10,   -21,     1,    -1,  
				  30,    -8,    27,     0,    -6,    44,  
				 -15,   -21,    -5,    10,    11,    19,  
				 -20,   -16,     8,   -11,   -20,    35,  
				 -12,   -11,     7,    37,    -7,    -7,  
				   3,    -6,   -11,   -14,   -16,   -13,  
				 -27,   -59,    -5,   -44,   -31,   -32,  
				 -28,    53,     4,   -33,   -25,   -37,  
				 -24,    30,    27,   -42,    29,   -31,  

				 -19,    61,    36,   -20,     6,    50,  
				 -27,    34,   -26,   -20,    90,     7,  
				 -30,    10,    14,    19,     3,   -26,  
				  47,    11,    33,    35,   -67,    -2,  
				 -28,    32,    -3,    10,   -15,    39,  
				 -19,   -32,    40,    22,    11,    27,  
				  -7,    38,   -11,    20,   -42,    32,  
				  12,   -20,     9,    13,    43,   -15,  
				   0,     1,    51,    -8,     8,   -17,  
				 -58,   -41,    -9,     1,    48,   -64,  
				 -29,    26,    48,   -19,    16,   -27,  
				 -21,   -28,    18,   -26,    36,   -13,  
				  14,    -7,    22,   -17,    13,    -7,  
				 -36,     8,    16,   -80,    -7,   -41,  
				   9,     5,    40,     2,   -61,   -50,  
				 -26,    20,    -5,   -17,    21,    36,  

				  45,    37,     0,   -14,   -20,    25,  
				  18,   -25,    -5,    24,    56,   -17,  
				 -19,    11,   -56,    -6,   -33,   -35,  
				  17,    -8,    19,    16,   -23,     0,  
				  -4,     6,   -43,    27,   -21,    21,  
				  44,   -32,    31,    -8,    10,    -1,  
				 -17,    30,    31,    25,   -12,   -11,  
				  -4,   -24,    22,   -27,    24,    11,  
				  18,   -30,    38,   -10,     0,    28,  
				   7,    -8,    12,    -9,    70,    -4,  
				 -20,   -21,    -8,     3,    18,     0,  
				 -32,   -25,   -24,    17,   -15,    -1,  
				  28,    -4,   -10,   -48,    82,   -33,  
				 -20,   -48,   -19,   -17,   -53,   -18,  
				  30,    22,    40,     6,   -22,    36,  
				   6,    16,   -29,    36,    20,     7
			};
	logic [0:27][0:27][0:5][31:0]	conv1 = {		
	 0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  

     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  

     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  

     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  

     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  

     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
    -7,       6,       4,       6,       0,      -7,  
   -17,      19,      19,      25,      -1,     -21,  
    -4,       8,      28,      50,      18,      -3,  
    17,     -21,      24,      73,      49,      26,  
    35,     -38,      25,      88,      44,      46,  
    38,     -42,      23,      84,      36,      67,  
    28,     -29,      17,      59,      14,      44,  
    16,     -15,      13,      36,       3,      36,  
     5,      -5,       5,      14,      -1,      11,  
     1,       0,       3,       5,      -2,       6,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  

     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
   -18,      24,      32,      17,     -12,     -21,  
   -12,      46,      97,      63,     -38,     -42,  
    54,      -5,     127,     140,       4,       4,  
   110,     -63,     155,     212,      18,      24,  
   132,     -86,     183,     254,      29,      63,  
   136,     -81,     174,     230,      34,      74,  
   105,     -75,     135,     198,      54,      79,  
    85,     -59,      99,     162,      53,      80,  
    51,     -44,      71,     147,      47,      70,  
    41,     -34,      58,     134,      44,      66,  
    33,     -34,      48,     130,      47,      60,  
    33,     -34,      48,     130,      47,      60,  
    33,     -34,      48,     130,      47,      60,  
    33,     -34,      48,     130,      47,      60,  
    36,     -36,      47,     128,      47,      63,  
    47,     -47,      37,     115,      47,      75,  
    48,     -53,      21,      91,      42,      79,  
    30,     -32,      16,      61,      11,      51,  
    12,      -8,      14,      33,      -6,      30,  
     2,       0,       4,       7,      -3,       8,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  

     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,      32,      68,      -3,     -46,     -15,  
    45,      50,     150,      35,    -106,     -35,  
   167,     -14,     206,     114,    -191,       7,  
   222,    -102,     253,     180,    -207,      42,  
   265,    -100,     307,     192,    -208,      80,  
   255,     -96,     324,     211,    -177,      87,  
   228,     -84,     302,     226,     -95,      79,  
   214,     -89,     292,     243,     -47,      77,  
   188,     -83,     273,     251,      -6,      66,  
   178,     -73,     268,     259,     -15,      56,  
   169,     -77,     258,     268,      -5,      61,  
   170,     -80,     255,     267,      -2,      57,  
   174,     -82,     256,     269,      -4,      64,  
   171,     -81,     255,     268,      -4,      62,  
   167,     -78,     251,     268,      -6,      55,  
   174,     -98,     211,     254,      18,      74,  
   166,    -116,     150,     201,      42,      99,  
   110,     -85,     101,     125,      33,      84,  
    53,     -23,      63,      56,      -7,      43,  
    14,       0,      21,      17,      -9,      22,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  

     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
    14,      48,      63,     -40,     -32,     -38,  
    83,      84,     127,     -82,     -95,     -42,  
   165,     -19,     145,     -71,    -222,     -49,  
   219,     -95,     160,     -49,    -286,      18,  
   273,    -104,     185,     -10,    -342,     117,  
   299,     -72,     212,      30,    -396,     156,  
   300,     -75,     230,      94,    -379,     161,  
   310,     -73,     267,     122,    -351,     154,  
   309,     -86,     300,     130,    -294,     143,  
   301,     -76,     331,     131,    -294,     105,  
   308,     -88,     337,     139,    -282,     108,  
   308,     -99,     331,     145,    -273,     103,  
   318,    -104,     333,     146,    -273,     116,  
   295,     -85,     343,     152,    -276,      97,  
   281,     -64,     362,     176,    -285,      75,  
   312,    -130,     306,     209,    -194,     145,  
   290,    -190,     208,     201,     -83,     161,  
   196,    -123,     166,     140,     -34,     156,  
    96,     -30,     117,      53,     -26,      88,  
    33,       2,      41,       5,     -15,      24,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  

     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
    10,      73,      54,     -72,      31,     -71,  
    36,      90,      86,    -167,      79,    -136,  
    66,     -27,      93,    -197,      39,    -150,  
    84,    -119,      35,    -147,      24,    -106,  
   119,     -52,      10,    -101,     -34,       1,  
   145,     -15,      20,     -94,    -110,      50,  
   180,     -18,      47,     -70,    -212,      71,  
   227,     -28,      65,     -57,    -277,     107,  
   252,     -34,      98,     -56,    -318,     114,  
   256,     -24,     133,     -74,    -315,     122,  
   280,     -46,     149,     -73,    -340,     104,  
   274,     -58,     144,     -60,    -332,     108,  
   275,     -55,     149,     -58,    -326,     107,  
   250,     -14,     210,     -44,    -353,      82,  
   277,     -18,     259,      18,    -346,      89,  
   377,    -157,     203,     133,    -319,     192,  
   348,    -248,     136,     215,    -244,     255,  
   243,    -124,     132,     152,    -166,     228,  
   123,      12,      94,      42,     -77,     158,  
    39,      16,      33,      -5,     -27,      39,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  

     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
    -8,      50,      27,     -56,      50,     -56,  
    12,      34,      69,    -112,     131,    -121,  
    -9,     -52,      24,    -128,     187,    -110,  
   -25,     -90,     -10,     -76,     197,    -107,  
   -11,     -19,     -23,     -76,     237,     -64,  
    -6,       9,     -10,    -110,     236,     -78,  
     7,     -13,      -2,    -129,     216,     -92,  
    29,     -35,     -21,    -115,     160,     -60,  
    51,     -34,     -10,    -106,     112,     -59,  
    73,      -1,     -11,    -117,     108,     -22,  
    84,     -17,       0,    -119,      64,     -31,  
    81,     -33,      -8,    -113,      71,     -32,  
    68,     -10,      19,     -84,      52,     -29,  
    78,      42,     131,     -57,       8,     -72,  
   211,      -5,     178,       8,       0,      19,  
   324,    -221,     107,     137,     -96,     118,  
   268,    -276,      44,     209,    -152,     235,  
   190,     -89,      60,     141,    -130,     264,  
   116,      63,      30,      38,     -67,     183,  
    28,      45,       3,       4,     -29,      59,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  

     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
    -3,      10,       4,     -12,      13,     -12,  
     0,       7,      18,     -28,      40,     -32,  
    -2,     -21,       8,     -26,      63,     -27,  
   -20,     -26,     -13,     -17,      78,     -24,  
   -19,      -4,      -2,     -20,     101,     -33,  
   -17,       4,       9,     -51,     144,     -45,  
   -21,     -12,      13,     -70,     185,     -78,  
   -30,     -49,     -14,     -60,     211,     -61,  
   -38,     -45,     -20,     -52,     215,     -58,  
   -27,     -23,     -26,     -48,     239,     -49,  
   -29,     -15,     -23,     -65,     231,     -42,  
   -40,     -35,     -18,     -42,     230,     -61,  
   -41,      13,      54,      -1,     165,     -59,  
    42,      73,     186,      15,     146,     -92,  
   217,     -32,     194,      43,     137,     -39,  
   261,    -281,     132,     106,      50,      77,  
   199,    -315,      57,     149,     -16,     179,  
   132,     -48,       0,     118,     -45,     263,  
    66,      83,     -13,      54,     -32,     159,  
    12,      52,      -8,       5,       0,      49,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  

     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       2,       1,      -3,       3,      -3,  
    -2,       7,       7,     -14,      17,     -15,  
     2,     -11,       7,      -9,      25,     -12,  
   -11,      -9,      -8,     -11,      36,      -9,  
    -6,      -4,       2,      -6,      42,     -20,  
   -11,       0,       2,     -13,      60,     -12,  
   -32,      16,      45,      19,      31,     -43,  
    10,      73,     162,      43,     -13,     -65,  
   163,      81,     256,      19,      -5,     -55,  
   301,    -140,     253,      38,      -3,     -52,  
   261,    -339,     156,      77,     -33,      71,  
   158,    -250,      57,     125,     -41,     188,  
    96,      16,     -18,      86,     -18,     200,  
    27,      90,     -20,      30,      -3,     103,  
     2,      25,      -2,       0,      12,      21,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  

     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
   -11,      15,      21,      10,      -9,     -12,  
    -7,      65,     121,      29,     -60,     -52,  
    98,     113,     250,      24,     -64,     -88,  
   262,     -13,     269,       4,     -34,     -85,  
   303,    -272,     216,      32,     -55,       7,  
   223,    -343,     105,      91,     -82,     132,  
   124,     -97,     -18,     102,     -54,     237,  
    54,      77,     -28,      57,     -22,     164,  
    12,      59,      -6,       5,      12,      61,  
     0,       3,       0,       0,       2,       2,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  

     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
   -14,      33,      52,      11,     -29,     -25,  
    25,     109,     187,      11,     -84,     -87,  
   180,      85,     267,     -15,     -59,     -86,  
   302,    -158,     243,      -5,     -23,     -68,  
   250,    -347,     137,      48,     -30,      61,  
   143,    -224,      33,      99,     -47,     196,  
    91,      15,     -33,      86,     -33,     193,  
    27,      93,     -32,      35,      -9,     110,  
     4,      26,      -4,       2,       4,      23,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  

     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
   -11,      10,       9,       9,      -1,     -11,  
   -11,      71,     107,      11,     -47,     -56,  
    78,     132,     236,     -18,     -41,    -103,  
   248,     -23,     249,     -25,     -18,     -95,  
   274,    -294,     170,      31,     -25,       7,  
   195,    -326,      85,     100,     -40,     127,  
   109,     -74,     -26,     100,     -10,     233,  
    34,      73,     -42,      62,      -3,     143,  
     3,      57,     -13,      10,      26,      53,  
     0,       8,       0,       0,       6,       7,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  

     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
    -6,       5,       4,       5,       0,      -6,  
   -21,      35,      53,      28,     -22,     -28,  
    19,     101,     182,      23,     -38,     -85,  
   171,      78,     264,     -11,       9,     -90,  
   286,    -172,     230,      16,       6,     -60,  
   228,    -362,     116,      88,     -30,      69,  
   129,    -198,      17,     117,     -33,     204,  
    83,      43,     -28,      81,     -23,     189,  
    18,      89,     -21,      21,       1,      94,  
     1,      13,      -1,       0,       8,      11,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  

     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
    -1,       1,       1,       1,       0,      -1,  
   -19,      24,      32,      19,     -11,     -21,  
    -4,      63,     131,      50,     -59,     -50,  
   113,      91,     247,      43,     -35,     -65,  
   271,     -39,     266,      27,      -6,     -74,  
   278,    -286,     196,      54,     -26,      25,  
   184,    -322,      89,      97,     -46,     124,  
   104,     -61,     -20,      99,     -21,     222,  
    42,      86,     -26,      51,     -16,     136,  
     6,      50,      -7,       3,      17,      43,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  

     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
   -18,      17,      16,      15,      -2,     -19,  
   -15,      56,     102,      43,     -49,     -42,  
    75,      69,     210,      68,     -51,     -40,  
   237,      25,     271,      48,     -58,     -52,  
   312,    -184,     260,      51,     -46,     -17,  
   253,    -336,     153,      61,     -61,      84,  
   134,    -196,      26,     100,     -50,     199,  
    78,      38,     -31,      78,     -27,     176,  
    18,      88,     -20,      19,       2,      91,  
     0,      11,       0,       0,       8,       9,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  

     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
    -3,       3,       2,       2,       0,      -3,  
   -19,      40,      69,      23,     -35,     -28,  
    25,      85,     187,      55,     -75,     -77,  
   196,      65,     275,      50,     -67,     -47,  
   304,    -117,     277,      33,     -46,     -62,  
   298,    -293,     210,      34,     -69,      37,  
   190,    -289,      81,      84,     -69,     161,  
    96,     -43,     -39,      86,     -27,     211,  
    36,      85,     -30,      52,     -14,     131,  
     6,      49,      -7,       2,      16,      42,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  

     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
    -2,       2,       1,       2,       0,      -2,  
   -19,      22,      25,      21,      -6,     -22,  
    -2,      73,     138,      36,     -65,     -53,  
   132,      88,     247,      35,     -64,     -40,  
   286,     -48,     262,      20,     -69,     -66,  
   301,    -237,     238,      14,     -59,      -2,  
   227,    -326,     125,      46,     -58,     114,  
   118,    -132,     -16,      80,     -43,     205,  
    57,      50,     -50,      76,     -13,     169,  
    14,      82,     -21,      19,       5,      82,  
     0,      11,       0,       0,       8,       9,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  

     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
   -11,      12,      15,      10,      -4,     -12,  
   -15,      50,      93,      38,     -44,     -38,  
    61,     102,     226,      44,     -49,     -87,  
   225,      42,     269,      20,     -25,     -75,  
   315,    -199,     265,      20,     -43,     -43,  
   253,    -334,     142,      34,     -26,      61,  
   154,    -206,      26,      84,     -48,     201,  
    68,      -3,     -62,      85,      -7,     202,  
    16,      83,     -40,      49,       0,     107,  
     4,      40,      -4,       0,      17,      35,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  

     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
    -5,       4,       3,       4,       0,      -5,  
   -19,      36,      56,      23,     -26,     -29,  
    20,      75,     167,      52,     -72,     -56,  
   159,      99,     289,      41,     -59,     -76,  
   303,     -96,     299,      53,     -23,     -82,  
   297,    -332,     202,      61,      20,      60,  
   201,    -330,      89,     121,       6,     155,  
   113,     -57,     -16,     118,      -8,     241,  
    31,      73,     -44,      71,      -3,     138,  
     4,      58,     -14,      10,      20,      52,  
     0,       6,       0,       0,       5,       5,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  

     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
   -10,      14,      21,       9,      -9,     -11,  
    -6,      66,     121,      26,     -58,     -54,  
    93,     111,     248,      34,     -77,     -86,  
   239,      29,     329,      31,     -84,    -103,  
   340,    -239,     306,      90,     -66,     -23,  
   331,    -407,     169,     163,     -41,     165,  
   181,    -207,      38,     185,     -19,     254,  
    96,      42,      15,     104,     -18,     211,  
    20,      72,      -4,      22,      13,      82,  
     1,      15,       0,       0,      11,      12,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  

     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
    -6,      25,      44,       3,     -27,     -17,  
    23,     108,     177,      -4,     -81,     -86,  
   152,     116,     290,     -20,     -87,    -123,  
   308,     -97,     347,      -9,     -90,    -105,  
   357,    -362,     220,      96,     -76,      84,  
   288,    -343,     108,     198,    -163,     215,  
   162,     -63,      33,     151,     -62,     273,  
    92,      92,      31,      31,     -36,     163,  
    18,      36,       7,      -1,       1,      39,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  

     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     9,      36,      57,     -25,     -29,     -25,  
    63,     126,     181,    -102,     -59,    -100,  
   181,      59,     261,    -134,    -104,    -162,  
   266,    -146,     247,    -106,    -120,    -134,  
   273,    -319,     111,      15,    -121,      71,  
   181,    -215,       8,      79,    -137,     209,  
   121,       1,     -29,      77,     -62,     225,  
    59,      98,      -9,      23,     -33,     155,  
     9,      23,       0,       1,      -5,      27,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  

     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     8,      50,      43,     -50,       8,     -48,  
    47,     118,     116,    -166,      34,    -131,  
   115,      12,     143,    -224,       1,    -157,  
   128,    -168,      56,    -178,      -8,     -92,  
   108,    -242,     -53,     -30,     -11,      66,  
    68,     -96,     -95,      51,     -12,     214,  
    49,      30,     -70,      89,     -22,     167,  
    22,      91,     -32,      28,      -3,      96,  
     3,      19,      -4,       2,       0,      17,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  

     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,      47,      29,     -49,      37,     -49,  
    13,      82,      76,    -146,     126,    -143,  
    13,      -9,      66,    -196,     181,    -174,  
    -3,    -157,     -18,    -106,     154,    -104,  
    12,    -152,     -83,      41,      89,      32,  
     3,     -10,    -123,      90,      63,     130,  
    -7,      69,     -63,      58,      26,      91,  
     0,      43,      -9,       7,      31,      40,  
     0,       7,       0,       0,       5,       6,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0,  
     0,       0,       0,       0,       0,       0 
		};
			
		
		go		 <= 0;
		en		 <= 0;
		first_data <= 0;
		last_data <= 0;
		data_i <= 0;
		weight <= 0;
		bias <= 0;
		@cb;
		@cb;
		@cb;
		@cb;
		
		for (int row = 0; row<32-4; row++) 
			for (int col = 0; col<32-4; col++) 
				for (int i = 0; i<5; i++) begin	
					for (int j = 0; j<5; j++) begin	
						en		 <= 1;
						if (i==0 && j ==0)
							first_data <= 1;
						else 
							first_data <= 0;
						if (i==4 && j ==4)
							last_data <= 1;
						else 
							last_data <= 0;
						data_i <= test[row + i][col +j];
						for(int w =0; w <`OUTPUT_NUM; w++ )
							weight[w] <= weight0[i][j][w];
						@cb;
					end
				end
		en		 <= 0;
	/*	
		go		 <= 0;
		en		 <= 0;
		first_data <= 0;
		last_data <= 0;
		data_i <= 0;
		weight <= 0;
		bias <= 0;
		@cb;
		@cb;
		go		 <= 1;
		@cb;
		go		 <= 0;
		@cb;
		
		for (int i = 0; i<9; i++) begin
			en		 <= 1;
			if(i == 0) first_data <= 1;
			else 		first_data <= 0;
			
			if(i == 8)  last_data <= 1;
			else 		last_data <= 0;
			
			for(int j = 0; j < `KERNEL_SIZE_SQ; j++) begin
				data_i[j] <= 1;
				weight[j] <= 1;
			end
			@cb;
		end
		en		 <= 0;
		last_data		 <= 0;
		first_data		 <= 0;
		
		@cb;
		@cb;
		@cb;
		@cb;
		@cb;
		@cb;
		@cb;
		@cb;
		@cb;
		@cb;
		@cb;
		@cb;
		@cb;
		@cb;
		@cb;
		@cb;
		go		 <= 1;
		@cb;
		go		 <= 0;
		@cb;
		for (int i = 0; i<3; i++) begin
			en		 <= 1;
			first_data <= 0;
			for(int j = 0; j < `KERNEL_SIZE_SQ; j++) begin
				data_i[j] <= 2;
				weight[j] <= 1;
			end
			@cb;
		end
		en		 <= 0;
		@cb;
		@cb;
		@cb;
		@cb;
		@cb;
		@cb;
		@cb;
		@cb;
		@cb;
		@cb;
		@cb;
		@cb;
		@cb;
		@cb;
		@cb;
		@cb;
		@cb;
		go		 <= 1;
		@cb;
		go		 <= 0;
		@cb;
		for (int i = 0; i<3; i++) begin
			en		 <= 1;
			first_data <= 0;
			if(i == 0)  last_data <= 1;
			else 		last_data <= 0;
			for(int j = 0; j < `KERNEL_SIZE_SQ; j++) begin
				data_i[j] <= 3;
				weight[j] <= 1;
			end
			@cb;
		end
			en		 <= 0;
		@cb;
		
		@cb;
		@cb;
		@cb;
		@cb;
		@cb;
		@cb;
		@cb;
		@cb;
		@cb;
		@cb;
		@cb;
		@cb;
		@cb;
		@cb;
		@cb;
		@cb;
		@cb;
	*/	
		

	endtask
	
	
endinterface
